<svg xmlns="http://www.w3.org/2000/svg" version="1.1" xmlns:xlink="http://www.w3.org/1999/xlink" xmlns:svgjs="http://svgjs.com/svgjs" width="2560" height="1440" preserveAspectRatio="none" viewBox="0 0 2560 1440"><g mask="url(&quot;#SvgjsMask1198&quot;)" fill="none"><rect width="2560" height="1440" x="0" y="0" fill="rgba(31, 32, 41, 1)"></rect><use xlink:href="#SvgjsSymbol1205" x="0" y="0"></use><use xlink:href="#SvgjsSymbol1205" x="0" y="720"></use><use xlink:href="#SvgjsSymbol1205" x="720" y="0"></use><use xlink:href="#SvgjsSymbol1205" x="720" y="720"></use><use xlink:href="#SvgjsSymbol1205" x="1440" y="0"></use><use xlink:href="#SvgjsSymbol1205" x="1440" y="720"></use><use xlink:href="#SvgjsSymbol1205" x="2160" y="0"></use><use xlink:href="#SvgjsSymbol1205" x="2160" y="720"></use></g><defs><mask id="SvgjsMask1198"><rect width="2560" height="1440" fill="#ffffff"></rect></mask><path d="M-1 0 a1 1 0 1 0 2 0 a1 1 0 1 0 -2 0z" id="SvgjsPath1204"></path><path d="M-3 0 a3 3 0 1 0 6 0 a3 3 0 1 0 -6 0z" id="SvgjsPath1199"></path><path d="M-5 0 a5 5 0 1 0 10 0 a5 5 0 1 0 -10 0z" id="SvgjsPath1202"></path><path d="M2 -2 L-2 2z" id="SvgjsPath1201"></path><path d="M6 -6 L-6 6z" id="SvgjsPath1200"></path><path d="M30 -30 L-30 30z" id="SvgjsPath1203"></path></defs><symbol id="SvgjsSymbol1205"><use xlink:href="#SvgjsPath1199" x="30" y="30" stroke="rgba(43, 44, 55, 1)"></use><use xlink:href="#SvgjsPath1200" x="30" y="90" stroke="rgba(43, 44, 55, 1)"></use><use xlink:href="#SvgjsPath1201" x="30" y="150" stroke="rgba(43, 44, 55, 1)"></use><use xlink:href="#SvgjsPath1200" x="30" y="210" stroke="rgba(43, 44, 55, 1)"></use><use xlink:href="#SvgjsPath1202" x="30" y="270" stroke="rgba(43, 44, 55, 1)"></use><use xlink:href="#SvgjsPath1202" x="30" y="330" stroke="rgba(43, 44, 55, 1)"></use><use xlink:href="#SvgjsPath1201" x="30" y="390" stroke="rgba(43, 44, 55, 1)"></use><use xlink:href="#SvgjsPath1199" x="30" y="450" stroke="rgba(43, 44, 55, 1)"></use><use xlink:href="#SvgjsPath1202" x="30" y="510" stroke="rgba(43, 44, 55, 1)"></use><use xlink:href="#SvgjsPath1199" x="30" y="570" stroke="rgba(43, 44, 55, 1)"></use><use xlink:href="#SvgjsPath1201" x="30" y="630" stroke="rgba(43, 44, 55, 1)"></use><use xlink:href="#SvgjsPath1201" x="30" y="690" stroke="rgba(43, 44, 55, 1)"></use><use xlink:href="#SvgjsPath1203" x="90" y="30" stroke="rgba(43, 44, 55, 1)" stroke-width="3"></use><use xlink:href="#SvgjsPath1204" x="90" y="90" stroke="rgba(43, 44, 55, 1)"></use><use xlink:href="#SvgjsPath1200" x="90" y="150" stroke="rgba(43, 44, 55, 1)"></use><use xlink:href="#SvgjsPath1201" x="90" y="210" stroke="rgba(43, 44, 55, 1)"></use><use xlink:href="#SvgjsPath1202" x="90" y="270" stroke="rgba(43, 44, 55, 1)"></use><use xlink:href="#SvgjsPath1200" x="90" y="330" stroke="rgba(43, 44, 55, 1)"></use><use xlink:href="#SvgjsPath1199" x="90" y="390" stroke="rgba(43, 44, 55, 1)"></use><use xlink:href="#SvgjsPath1202" x="90" y="450" stroke="rgba(43, 44, 55, 1)"></use><use xlink:href="#SvgjsPath1203" x="90" y="510" stroke="rgba(43, 44, 55, 1)" stroke-width="3"></use><use xlink:href="#SvgjsPath1200" x="90" y="570" stroke="rgba(43, 44, 55, 1)"></use><use xlink:href="#SvgjsPath1200" x="90" y="630" stroke="rgba(43, 44, 55, 1)"></use><use xlink:href="#SvgjsPath1201" x="90" y="690" stroke="rgba(43, 44, 55, 1)"></use><use xlink:href="#SvgjsPath1204" x="150" y="30" stroke="rgba(43, 44, 55, 1)"></use><use xlink:href="#SvgjsPath1202" x="150" y="90" stroke="rgba(43, 44, 55, 1)"></use><use xlink:href="#SvgjsPath1200" x="150" y="150" stroke="rgba(43, 44, 55, 1)"></use><use xlink:href="#SvgjsPath1200" x="150" y="210" stroke="rgba(43, 44, 55, 1)"></use><use xlink:href="#SvgjsPath1200" x="150" y="270" stroke="rgba(43, 44, 55, 1)"></use><use xlink:href="#SvgjsPath1202" x="150" y="330" stroke="rgba(43, 44, 55, 1)"></use><use xlink:href="#SvgjsPath1202" x="150" y="390" stroke="rgba(43, 44, 55, 1)"></use><use xlink:href="#SvgjsPath1204" x="150" y="450" stroke="rgba(43, 44, 55, 1)"></use><use xlink:href="#SvgjsPath1202" x="150" y="510" stroke="rgba(43, 44, 55, 1)"></use><use xlink:href="#SvgjsPath1204" x="150" y="570" stroke="rgba(43, 44, 55, 1)"></use><use xlink:href="#SvgjsPath1202" x="150" y="630" stroke="rgba(43, 44, 55, 1)"></use><use xlink:href="#SvgjsPath1204" x="150" y="690" stroke="rgba(43, 44, 55, 1)"></use><use xlink:href="#SvgjsPath1199" x="210" y="30" stroke="rgba(43, 44, 55, 1)"></use><use xlink:href="#SvgjsPath1200" x="210" y="90" stroke="rgba(43, 44, 55, 1)"></use><use xlink:href="#SvgjsPath1200" x="210" y="150" stroke="rgba(43, 44, 55, 1)"></use><use xlink:href="#SvgjsPath1203" x="210" y="210" stroke="rgba(43, 44, 55, 1)" stroke-width="3"></use><use xlink:href="#SvgjsPath1200" x="210" y="270" stroke="rgba(43, 44, 55, 1)"></use><use xlink:href="#SvgjsPath1202" x="210" y="330" stroke="rgba(43, 44, 55, 1)"></use><use xlink:href="#SvgjsPath1200" x="210" y="390" stroke="rgba(43, 44, 55, 1)"></use><use xlink:href="#SvgjsPath1199" x="210" y="450" stroke="rgba(43, 44, 55, 1)"></use><use xlink:href="#SvgjsPath1204" x="210" y="510" stroke="rgba(43, 44, 55, 1)"></use><use xlink:href="#SvgjsPath1204" x="210" y="570" stroke="rgba(43, 44, 55, 1)"></use><use xlink:href="#SvgjsPath1200" x="210" y="630" stroke="rgba(43, 44, 55, 1)"></use><use xlink:href="#SvgjsPath1200" x="210" y="690" stroke="rgba(43, 44, 55, 1)"></use><use xlink:href="#SvgjsPath1201" x="270" y="30" stroke="rgba(43, 44, 55, 1)"></use><use xlink:href="#SvgjsPath1203" x="270" y="90" stroke="rgba(43, 44, 55, 1)" stroke-width="3"></use><use xlink:href="#SvgjsPath1202" x="270" y="150" stroke="rgba(43, 44, 55, 1)"></use><use xlink:href="#SvgjsPath1201" x="270" y="210" stroke="rgba(43, 44, 55, 1)"></use><use xlink:href="#SvgjsPath1200" x="270" y="270" stroke="rgba(43, 44, 55, 1)"></use><use xlink:href="#SvgjsPath1202" x="270" y="330" stroke="rgba(43, 44, 55, 1)"></use><use xlink:href="#SvgjsPath1201" x="270" y="390" stroke="rgba(43, 44, 55, 1)"></use><use xlink:href="#SvgjsPath1200" x="270" y="450" stroke="rgba(43, 44, 55, 1)"></use><use xlink:href="#SvgjsPath1200" x="270" y="510" stroke="rgba(43, 44, 55, 1)"></use><use xlink:href="#SvgjsPath1202" x="270" y="570" stroke="rgba(43, 44, 55, 1)"></use><use xlink:href="#SvgjsPath1200" x="270" y="630" stroke="rgba(43, 44, 55, 1)"></use><use xlink:href="#SvgjsPath1200" x="270" y="690" stroke="rgba(43, 44, 55, 1)"></use><use xlink:href="#SvgjsPath1201" x="330" y="30" stroke="rgba(43, 44, 55, 1)"></use><use xlink:href="#SvgjsPath1200" x="330" y="90" stroke="rgba(43, 44, 55, 1)"></use><use xlink:href="#SvgjsPath1200" x="330" y="150" stroke="rgba(43, 44, 55, 1)"></use><use xlink:href="#SvgjsPath1201" x="330" y="210" stroke="rgba(43, 44, 55, 1)"></use><use xlink:href="#SvgjsPath1202" x="330" y="270" stroke="rgba(43, 44, 55, 1)"></use><use xlink:href="#SvgjsPath1201" x="330" y="330" stroke="rgba(43, 44, 55, 1)"></use><use xlink:href="#SvgjsPath1200" x="330" y="390" stroke="rgba(43, 44, 55, 1)"></use><use xlink:href="#SvgjsPath1202" x="330" y="450" stroke="rgba(43, 44, 55, 1)"></use><use xlink:href="#SvgjsPath1202" x="330" y="510" stroke="rgba(43, 44, 55, 1)"></use><use xlink:href="#SvgjsPath1199" x="330" y="570" stroke="rgba(43, 44, 55, 1)"></use><use xlink:href="#SvgjsPath1200" x="330" y="630" stroke="rgba(43, 44, 55, 1)"></use><use xlink:href="#SvgjsPath1200" x="330" y="690" stroke="rgba(43, 44, 55, 1)"></use><use xlink:href="#SvgjsPath1202" x="390" y="30" stroke="rgba(43, 44, 55, 1)"></use><use xlink:href="#SvgjsPath1199" x="390" y="90" stroke="rgba(43, 44, 55, 1)"></use><use xlink:href="#SvgjsPath1203" x="390" y="150" stroke="rgba(43, 44, 55, 1)" stroke-width="3"></use><use xlink:href="#SvgjsPath1201" x="390" y="210" stroke="rgba(43, 44, 55, 1)"></use><use xlink:href="#SvgjsPath1202" x="390" y="270" stroke="rgba(43, 44, 55, 1)"></use><use xlink:href="#SvgjsPath1202" x="390" y="330" stroke="rgba(43, 44, 55, 1)"></use><use xlink:href="#SvgjsPath1203" x="390" y="390" stroke="rgba(43, 44, 55, 1)" stroke-width="3"></use><use xlink:href="#SvgjsPath1200" x="390" y="450" stroke="rgba(43, 44, 55, 1)"></use><use xlink:href="#SvgjsPath1201" x="390" y="510" stroke="rgba(43, 44, 55, 1)"></use><use xlink:href="#SvgjsPath1204" x="390" y="570" stroke="rgba(43, 44, 55, 1)"></use><use xlink:href="#SvgjsPath1201" x="390" y="630" stroke="rgba(43, 44, 55, 1)"></use><use xlink:href="#SvgjsPath1204" x="390" y="690" stroke="rgba(43, 44, 55, 1)"></use><use xlink:href="#SvgjsPath1200" x="450" y="30" stroke="rgba(43, 44, 55, 1)"></use><use xlink:href="#SvgjsPath1204" x="450" y="90" stroke="rgba(43, 44, 55, 1)"></use><use xlink:href="#SvgjsPath1201" x="450" y="150" stroke="rgba(43, 44, 55, 1)"></use><use xlink:href="#SvgjsPath1199" x="450" y="210" stroke="rgba(43, 44, 55, 1)"></use><use xlink:href="#SvgjsPath1203" x="450" y="270" stroke="rgba(43, 44, 55, 1)" stroke-width="3"></use><use xlink:href="#SvgjsPath1202" x="450" y="330" stroke="rgba(43, 44, 55, 1)"></use><use xlink:href="#SvgjsPath1202" x="450" y="390" stroke="rgba(43, 44, 55, 1)"></use><use xlink:href="#SvgjsPath1202" x="450" y="450" stroke="rgba(43, 44, 55, 1)"></use><use xlink:href="#SvgjsPath1202" x="450" y="510" stroke="rgba(43, 44, 55, 1)"></use><use xlink:href="#SvgjsPath1203" x="450" y="570" stroke="rgba(43, 44, 55, 1)" stroke-width="3"></use><use xlink:href="#SvgjsPath1200" x="450" y="630" stroke="rgba(43, 44, 55, 1)"></use><use xlink:href="#SvgjsPath1200" x="450" y="690" stroke="rgba(43, 44, 55, 1)"></use><use xlink:href="#SvgjsPath1200" x="510" y="30" stroke="rgba(43, 44, 55, 1)"></use><use xlink:href="#SvgjsPath1201" x="510" y="90" stroke="rgba(43, 44, 55, 1)"></use><use xlink:href="#SvgjsPath1201" x="510" y="150" stroke="rgba(43, 44, 55, 1)"></use><use xlink:href="#SvgjsPath1200" x="510" y="210" stroke="rgba(43, 44, 55, 1)"></use><use xlink:href="#SvgjsPath1199" x="510" y="270" stroke="rgba(43, 44, 55, 1)"></use><use xlink:href="#SvgjsPath1202" x="510" y="330" stroke="rgba(43, 44, 55, 1)"></use><use xlink:href="#SvgjsPath1202" x="510" y="390" stroke="rgba(43, 44, 55, 1)"></use><use xlink:href="#SvgjsPath1199" x="510" y="450" stroke="rgba(43, 44, 55, 1)"></use><use xlink:href="#SvgjsPath1202" x="510" y="510" stroke="rgba(43, 44, 55, 1)"></use><use xlink:href="#SvgjsPath1204" x="510" y="570" stroke="rgba(43, 44, 55, 1)"></use><use xlink:href="#SvgjsPath1202" x="510" y="630" stroke="rgba(43, 44, 55, 1)"></use><use xlink:href="#SvgjsPath1202" x="510" y="690" stroke="rgba(43, 44, 55, 1)"></use><use xlink:href="#SvgjsPath1202" x="570" y="30" stroke="rgba(43, 44, 55, 1)"></use><use xlink:href="#SvgjsPath1202" x="570" y="90" stroke="rgba(43, 44, 55, 1)"></use><use xlink:href="#SvgjsPath1201" x="570" y="150" stroke="rgba(43, 44, 55, 1)"></use><use xlink:href="#SvgjsPath1200" x="570" y="210" stroke="rgba(43, 44, 55, 1)"></use><use xlink:href="#SvgjsPath1204" x="570" y="270" stroke="rgba(43, 44, 55, 1)"></use><use xlink:href="#SvgjsPath1202" x="570" y="330" stroke="rgba(43, 44, 55, 1)"></use><use xlink:href="#SvgjsPath1201" x="570" y="390" stroke="rgba(43, 44, 55, 1)"></use><use xlink:href="#SvgjsPath1201" x="570" y="450" stroke="rgba(43, 44, 55, 1)"></use><use xlink:href="#SvgjsPath1201" x="570" y="510" stroke="rgba(43, 44, 55, 1)"></use><use xlink:href="#SvgjsPath1202" x="570" y="570" stroke="rgba(43, 44, 55, 1)"></use><use xlink:href="#SvgjsPath1200" x="570" y="630" stroke="rgba(43, 44, 55, 1)"></use><use xlink:href="#SvgjsPath1200" x="570" y="690" stroke="rgba(43, 44, 55, 1)"></use><use xlink:href="#SvgjsPath1202" x="630" y="30" stroke="rgba(43, 44, 55, 1)"></use><use xlink:href="#SvgjsPath1200" x="630" y="90" stroke="rgba(43, 44, 55, 1)"></use><use xlink:href="#SvgjsPath1200" x="630" y="150" stroke="rgba(43, 44, 55, 1)"></use><use xlink:href="#SvgjsPath1200" x="630" y="210" stroke="rgba(43, 44, 55, 1)"></use><use xlink:href="#SvgjsPath1204" x="630" y="270" stroke="rgba(43, 44, 55, 1)"></use><use xlink:href="#SvgjsPath1200" x="630" y="330" stroke="rgba(43, 44, 55, 1)"></use><use xlink:href="#SvgjsPath1204" x="630" y="390" stroke="rgba(43, 44, 55, 1)"></use><use xlink:href="#SvgjsPath1202" x="630" y="450" stroke="rgba(43, 44, 55, 1)"></use><use xlink:href="#SvgjsPath1202" x="630" y="510" stroke="rgba(43, 44, 55, 1)"></use><use xlink:href="#SvgjsPath1200" x="630" y="570" stroke="rgba(43, 44, 55, 1)"></use><use xlink:href="#SvgjsPath1203" x="630" y="630" stroke="rgba(43, 44, 55, 1)" stroke-width="3"></use><use xlink:href="#SvgjsPath1199" x="630" y="690" stroke="rgba(43, 44, 55, 1)"></use><use xlink:href="#SvgjsPath1202" x="690" y="30" stroke="rgba(43, 44, 55, 1)"></use><use xlink:href="#SvgjsPath1202" x="690" y="90" stroke="rgba(43, 44, 55, 1)"></use><use xlink:href="#SvgjsPath1204" x="690" y="150" stroke="rgba(43, 44, 55, 1)"></use><use xlink:href="#SvgjsPath1202" x="690" y="210" stroke="rgba(43, 44, 55, 1)"></use><use xlink:href="#SvgjsPath1202" x="690" y="270" stroke="rgba(43, 44, 55, 1)"></use><use xlink:href="#SvgjsPath1200" x="690" y="330" stroke="rgba(43, 44, 55, 1)"></use><use xlink:href="#SvgjsPath1200" x="690" y="390" stroke="rgba(43, 44, 55, 1)"></use><use xlink:href="#SvgjsPath1200" x="690" y="450" stroke="rgba(43, 44, 55, 1)"></use><use xlink:href="#SvgjsPath1199" x="690" y="510" stroke="rgba(43, 44, 55, 1)"></use><use xlink:href="#SvgjsPath1201" x="690" y="570" stroke="rgba(43, 44, 55, 1)"></use><use xlink:href="#SvgjsPath1200" x="690" y="630" stroke="rgba(43, 44, 55, 1)"></use><use xlink:href="#SvgjsPath1202" x="690" y="690" stroke="rgba(43, 44, 55, 1)"></use></symbol></svg>
